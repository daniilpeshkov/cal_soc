//------------------------------------------------------
//	Wishbone rom
//------------------------------------------------------
//	author:  	Peshkov Daniil
//	email:  	daniil.peshkov@spbpu.com
//------------------------------------------------------


module moduleName #(
    parameters
) (
    ports
);
    
endmodule
