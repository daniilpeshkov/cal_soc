
module tb_ch_measure_ctl();




endmodule